`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/01/26 17:06:49
// Design Name: 
// Module Name: ifm_controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ifm_controller(
    input clk,
    input rst_n,
    input is_conv_3,
    input is_maxpooling,
    input [10:0] ifm_channel,
    input [10:0] ofm_channel,
    input [8:0] ifm_width,
    
    input          temp_valid,
    output         temp_hs,
    input [15:0]   temp_data_0, temp_data_1, temp_data_2, temp_data_3, 
                   temp_data_4, temp_data_5, temp_data_6, temp_data_7, 
                   temp_data_8, temp_data_9, temp_data_10, temp_data_11, 
                   temp_data_12, temp_data_13, temp_data_14, temp_data_15,
                   temp_data_16, temp_data_17, temp_data_18, temp_data_19,
                   temp_data_20, temp_data_21, temp_data_22, temp_data_23, 
                   temp_data_24, temp_data_25, temp_data_26, temp_data_27, 
                   temp_data_28, temp_data_29, temp_data_30, temp_data_31,
                   temp_data_32, temp_data_33, temp_data_34, temp_data_35,
                   temp_data_36, temp_data_37, temp_data_38, temp_data_39,
                   temp_data_40, temp_data_41, temp_data_42, temp_data_43,
    
    output reg        conv3_ifm_valid,               
    input             conv3_ifm_weight_hs,
    output reg [15:0]  ifm_data_0,  ifm_data_1,  ifm_data_2,  ifm_data_3,  ifm_data_4,  ifm_data_5,  ifm_data_6,  ifm_data_7,  ifm_data_8,  ifm_data_9, ifm_data_10,  ifm_data_11, ifm_data_12, ifm_data_13, ifm_data_14,
                       ifm_data_15, ifm_data_16, ifm_data_17, ifm_data_18, ifm_data_19, ifm_data_20, ifm_data_21, ifm_data_22, ifm_data_23, ifm_data_24, ifm_data_25, ifm_data_26, ifm_data_27, ifm_data_28, ifm_data_29,
                       ifm_data_30, ifm_data_31, ifm_data_32, ifm_data_33, ifm_data_34, ifm_data_35, ifm_data_36, ifm_data_37, ifm_data_38, ifm_data_39, ifm_data_40, ifm_data_41, ifm_data_42, ifm_data_43, ifm_data_44
    );
    
    
    reg last_col_2cycle;
    reg last_col_2cycle_buf;
    wire last_col;
    wire conv3_row1;
    wire conv3_reuse;
    wire conv3_rowlast;
    reg buf_conv3_rowlast;
    wire [4:0] w_cnt;
    wire [1:0] remain;
    wire [1:0] remain_13;
    wire [4:0] w_finish_cnt;
    wire temp_ready = (conv3_ifm_valid ==0 ||conv3_ifm_weight_hs)&(conv3_row1||conv3_reuse &!(last_col_2cycle||last_col_2cycle_buf));
    
    reg bram_hs;
    
    ifm_remain_controller ifm_remain_controller(
    .clk(clk),
    .rst_n(rst_n),
    .is_conv_3(is_conv_3),
    .last_col(last_col),
    .conv3_row1(conv3_row1),
    .conv3_reuse(conv3_reuse),
    .conv3_rowlast(conv3_rowlast),
    .w_cnt(w_cnt),
    .remain(remain),
    .remain_13(remain_13),
    .w_finish_cnt(w_finish_cnt),
    .temp_hs(temp_hs),
    .ifm_width(ifm_width),
    .ifm_channel(ifm_channel),
    .ofm_channel(ofm_channel),
    .bram_hs(bram_hs)
    );

    reg read_flag;
    reg buf_read_flag;

    
    wire [23:0] reuse_data_2bram [0:19];
    wire [23:0] reuse_data_2ifm0 [0:19];
    wire [23:0] reuse_data_2ifm1 [0:19];
    
    assign reuse_data_2bram[0] = {ifm_data_16[7:0],ifm_data_15}; assign reuse_data_2bram[1] = {ifm_data_17,ifm_data_16[15:8]};
    assign reuse_data_2bram[2] = {ifm_data_19[7:0],ifm_data_18}; assign reuse_data_2bram[3] = {ifm_data_20,ifm_data_19[15:8]};
    assign reuse_data_2bram[4] = {ifm_data_22[7:0],ifm_data_21}; assign reuse_data_2bram[5] = {ifm_data_23,ifm_data_22[15:8]};
    assign reuse_data_2bram[6] = {ifm_data_25[7:0],ifm_data_24}; assign reuse_data_2bram[7] = {ifm_data_26,ifm_data_25[15:8]};
    assign reuse_data_2bram[8] = {ifm_data_28[7:0],ifm_data_27}; assign reuse_data_2bram[9] = {ifm_data_29,ifm_data_28[15:8]};
    assign reuse_data_2bram[10] = {ifm_data_31[7:0],ifm_data_30}; assign reuse_data_2bram[11] = {ifm_data_32,ifm_data_31[15:8]};
    assign reuse_data_2bram[12] = {ifm_data_34[7:0],ifm_data_33}; assign reuse_data_2bram[13] = {ifm_data_35,ifm_data_34[15:8]};
    assign reuse_data_2bram[14] = {ifm_data_37[7:0],ifm_data_36}; assign reuse_data_2bram[15] = {ifm_data_38,ifm_data_37[15:8]};
    assign reuse_data_2bram[16] = {ifm_data_40[7:0],ifm_data_39}; assign reuse_data_2bram[17] = {ifm_data_41,ifm_data_40[15:8]};
    assign reuse_data_2bram[18] = {ifm_data_43[7:0],ifm_data_42}; assign reuse_data_2bram[19] = {ifm_data_44,ifm_data_43[15:8]};
    
    genvar i;
    generate
        for(i =0; i<20; i=i+1)begin:IFM_BRAM_0
             reuse_bram_controller#(.r_flag(1'b0))Reuse_BRAM_0_Controller
            (
            .clk(clk),
            .rst_n(rst_n),
            .read_flag(buf_read_flag),
            .bram_hs(bram_hs),
            .din(reuse_data_2bram[i]),
            .dout(reuse_data_2ifm0[i]),
            .conv3_reuse(conv3_reuse),
            .conv3_rowlast(conv3_rowlast),
            .temp_hs(temp_hs),
            .buf_conv3_rowlast(buf_conv3_rowlast)
            );
        end
    endgenerate
    //
    generate
        for(i =0; i<20; i=i+1)begin:IFM_BRAM_1
             reuse_bram_controller#(.r_flag(1'b1))Reuse_BRAM_1_Controller
            (
            .clk(clk),
            .rst_n(rst_n),
            .read_flag(buf_read_flag),
            .bram_hs(bram_hs),
            .din(reuse_data_2bram[i]),
            .dout(reuse_data_2ifm1[i]),
            .conv3_reuse(conv3_reuse),
            .conv3_rowlast(conv3_rowlast),
            .temp_hs(temp_hs),
            .buf_conv3_rowlast(buf_conv3_rowlast)
            );
        end
    endgenerate
    
    reg [1:0] low_last_ready_cnt;
    reg bram_temp_hs;
    
    assign temp_hs = temp_valid & temp_ready;
    
    always@(posedge clk)begin
        if(!rst_n)begin
            bram_temp_hs<=0;
            buf_conv3_rowlast <= 0;
            low_last_ready_cnt<=0;
            bram_hs<=0;
            read_flag <=0;
            buf_read_flag <=0;
            last_col_2cycle <=0;
            last_col_2cycle_buf <=0;
            conv3_ifm_valid <= 0;
            ifm_data_0<= 0; ifm_data_1<=0; ifm_data_2<=0;  ifm_data_3<=0;  ifm_data_4<=0;  ifm_data_5<=0;  ifm_data_6<=0;  ifm_data_7<=0;  ifm_data_8<=0; ifm_data_9<=0; ifm_data_10<=0; ifm_data_11<=0; ifm_data_12<=0; ifm_data_13<=0; ifm_data_14<=0;
            ifm_data_15<=0;  ifm_data_16<=0; ifm_data_17<=0;  ifm_data_18<=0;  ifm_data_19<=0;  ifm_data_20<=0;  ifm_data_21<=0;  ifm_data_22<=0;  ifm_data_23<=0; ifm_data_24<=0; ifm_data_25<=0; ifm_data_26<=0; ifm_data_27<=0; ifm_data_28<=0; ifm_data_29<=0;
            ifm_data_30<=0;  ifm_data_31<=0; ifm_data_32<=0;  ifm_data_33<=0;  ifm_data_34<=0;  ifm_data_35<=0;  ifm_data_36<=0;  ifm_data_37<=0;  ifm_data_38<=0; ifm_data_39<=0; ifm_data_40<=0; ifm_data_41<=0; ifm_data_42<=0; ifm_data_43<=0; ifm_data_44<=0;
        end else begin
            buf_conv3_rowlast <= conv3_rowlast;
            buf_read_flag <= read_flag;
            if(temp_hs)conv3_ifm_valid <=1;
            else if(conv3_ifm_weight_hs)conv3_ifm_valid <=0;
            else if(conv3_ifm_valid ==0 & buf_conv3_rowlast & bram_hs)conv3_ifm_valid <=1;
            
            if(conv3_rowlast & low_last_ready_cnt != 2) low_last_ready_cnt <= low_last_ready_cnt+1;//wrong
            else if (!conv3_rowlast) low_last_ready_cnt <= 0;
            
            if(conv3_rowlast & (low_last_ready_cnt < 2) & conv3_ifm_weight_hs) bram_temp_hs <=1;
            else if(low_last_ready_cnt ==2)bram_temp_hs <=0;

            if(temp_hs || (conv3_rowlast& (bram_temp_hs||conv3_ifm_weight_hs)& low_last_ready_cnt ==2))bram_hs<=1;
            else bram_hs<=0;
            
            if(last_col & temp_hs)begin
                last_col_2cycle<=1;
                read_flag <= read_flag+1;
            end else begin
                last_col_2cycle<=0;
            end
            last_col_2cycle_buf<=last_col_2cycle;
            
            if(conv3_row1 & temp_hs)begin
                ifm_data_0<= 1; ifm_data_1<=1; ifm_data_2<=1;  ifm_data_3<=1;  ifm_data_4<=1;  ifm_data_5<=1;  ifm_data_6<=1;  ifm_data_7<=1;  ifm_data_8<=1; ifm_data_9<=1; ifm_data_10<=1; ifm_data_11<=1; ifm_data_12<=1; ifm_data_13<=1; ifm_data_14<=1;
                case(ifm_width)
                    default:begin
                        if(w_cnt ==0)begin
                            ifm_data_15<=1;
                            ifm_data_30<=1;
                            ifm_data_16<=temp_data_0; ifm_data_17<=temp_data_1;  ifm_data_18<=temp_data_2;  ifm_data_19<=temp_data_3;  ifm_data_20<=temp_data_4;  ifm_data_21<=temp_data_5;  ifm_data_22<=temp_data_6;  ifm_data_23<=temp_data_7; ifm_data_24<=temp_data_8; ifm_data_25<=temp_data_9; ifm_data_26<=temp_data_10; ifm_data_27<=temp_data_11; ifm_data_28<=temp_data_12; ifm_data_29<=temp_data_13;
                            ifm_data_31<=temp_data_16; ifm_data_32<=temp_data_17;  ifm_data_33<=temp_data_18;  ifm_data_34<=temp_data_19;  ifm_data_35<=temp_data_20;  ifm_data_36<=temp_data_21;  ifm_data_37<=temp_data_22;  ifm_data_38<=temp_data_23; ifm_data_39<=temp_data_24; ifm_data_40<=temp_data_25; ifm_data_41<=temp_data_26; ifm_data_42<=temp_data_27; ifm_data_43<=temp_data_28; ifm_data_44<=temp_data_29;
                        end else if(w_cnt == w_finish_cnt)begin
                            ifm_data_29<=1;
                            ifm_data_44<=1;
                            ifm_data_15<=temp_data_2;  ifm_data_16<=temp_data_3; ifm_data_17<=temp_data_4;  ifm_data_18<=temp_data_5;  ifm_data_19<=temp_data_6;  ifm_data_20<=temp_data_7;  ifm_data_21<=temp_data_8;  ifm_data_22<=temp_data_9;  ifm_data_23<=temp_data_10; ifm_data_24<=temp_data_11; ifm_data_25<=temp_data_12; ifm_data_26<=temp_data_13; ifm_data_27<=temp_data_14; ifm_data_28<=temp_data_15;
                            ifm_data_30<=temp_data_18;  ifm_data_31<=temp_data_19; ifm_data_32<=temp_data_20;  ifm_data_33<=temp_data_21;  ifm_data_34<=temp_data_22;  ifm_data_35<=temp_data_23;  ifm_data_36<=temp_data_24;  ifm_data_37<=temp_data_25;  ifm_data_38<=temp_data_26; ifm_data_39<=temp_data_27; ifm_data_40<=temp_data_28; ifm_data_41<=temp_data_29; ifm_data_42<=temp_data_30; ifm_data_43<=temp_data_31;
                        end else begin
                            case(remain)
                                0:begin
                                    ifm_data_15<=temp_data_1;  ifm_data_16<=temp_data_2; ifm_data_17<=temp_data_3;  ifm_data_18<=temp_data_4;  ifm_data_19<=temp_data_5;  ifm_data_20<=temp_data_6;  ifm_data_21<=temp_data_7;  ifm_data_22<=temp_data_8;  ifm_data_23<=temp_data_9; ifm_data_24<=temp_data_10; ifm_data_25<=temp_data_11; ifm_data_26<=temp_data_12; ifm_data_27<=temp_data_13; ifm_data_28<=temp_data_14; ifm_data_29<=temp_data_15;
                                    ifm_data_30<=temp_data_17;  ifm_data_31<=temp_data_18; ifm_data_32<=temp_data_19;  ifm_data_33<=temp_data_20;  ifm_data_34<=temp_data_21;  ifm_data_35<=temp_data_22;  ifm_data_36<=temp_data_23;  ifm_data_37<=temp_data_24;  ifm_data_38<=temp_data_25; ifm_data_39<=temp_data_26; ifm_data_40<=temp_data_27; ifm_data_41<=temp_data_28; ifm_data_42<=temp_data_29; ifm_data_43<=temp_data_30; ifm_data_44<=temp_data_31;
                                end
                                1:begin
                                    ifm_data_15<=temp_data_0;  ifm_data_16<=temp_data_1; ifm_data_17<=temp_data_2;  ifm_data_18<=temp_data_3;  ifm_data_19<=temp_data_4;  ifm_data_20<=temp_data_5;  ifm_data_21<=temp_data_6;  ifm_data_22<=temp_data_7;  ifm_data_23<=temp_data_8; ifm_data_24<=temp_data_9; ifm_data_25<=temp_data_10; ifm_data_26<=temp_data_11; ifm_data_27<=temp_data_12; ifm_data_28<=temp_data_13; ifm_data_29<=temp_data_14;
                                    ifm_data_30<=temp_data_16;  ifm_data_31<=temp_data_17; ifm_data_32<=temp_data_18;  ifm_data_33<=temp_data_19;  ifm_data_34<=temp_data_20;  ifm_data_35<=temp_data_21;  ifm_data_36<=temp_data_22;  ifm_data_37<=temp_data_23;  ifm_data_38<=temp_data_24; ifm_data_39<=temp_data_25; ifm_data_40<=temp_data_26; ifm_data_41<=temp_data_27; ifm_data_42<=temp_data_28; ifm_data_43<=temp_data_29; ifm_data_44<=temp_data_30;
                                end
                                2:begin
                                    ifm_data_15<=temp_data_3;  ifm_data_16<=temp_data_4; ifm_data_17<=temp_data_5;  ifm_data_18<=temp_data_6;  ifm_data_19<=temp_data_7;  ifm_data_20<=temp_data_8;  ifm_data_21<=temp_data_9;  ifm_data_22<=temp_data_10;  ifm_data_23<=temp_data_11; ifm_data_24<=temp_data_12; ifm_data_25<=temp_data_13; ifm_data_26<=temp_data_14; ifm_data_27<=temp_data_15; ifm_data_28<=temp_data_16; ifm_data_29<=temp_data_17;
                                    ifm_data_30<=temp_data_23;  ifm_data_31<=temp_data_24; ifm_data_32<=temp_data_25;  ifm_data_33<=temp_data_26;  ifm_data_34<=temp_data_27;  ifm_data_35<=temp_data_28;  ifm_data_36<=temp_data_29;  ifm_data_37<=temp_data_30;  ifm_data_38<=temp_data_31; ifm_data_39<=temp_data_32; ifm_data_40<=temp_data_33; ifm_data_41<=temp_data_34; ifm_data_42<=temp_data_35; ifm_data_43<=temp_data_36; ifm_data_44<=temp_data_37;
                                end
                                3:begin
                                    ifm_data_15<=temp_data_2;  ifm_data_16<=temp_data_3; ifm_data_17<=temp_data_4;  ifm_data_18<=temp_data_5;  ifm_data_19<=temp_data_6;  ifm_data_20<=temp_data_7;  ifm_data_21<=temp_data_8;  ifm_data_22<=temp_data_9;  ifm_data_23<=temp_data_10; ifm_data_24<=temp_data_11; ifm_data_25<=temp_data_12; ifm_data_26<=temp_data_13; ifm_data_27<=temp_data_14; ifm_data_28<=temp_data_15; ifm_data_29<=temp_data_16;
                                    ifm_data_30<=temp_data_22;  ifm_data_31<=temp_data_23; ifm_data_32<=temp_data_24;  ifm_data_33<=temp_data_25;  ifm_data_34<=temp_data_26;  ifm_data_35<=temp_data_27;  ifm_data_36<=temp_data_28;  ifm_data_37<=temp_data_29;  ifm_data_38<=temp_data_30; ifm_data_39<=temp_data_31; ifm_data_40<=temp_data_32; ifm_data_41<=temp_data_33; ifm_data_42<=temp_data_34; ifm_data_43<=temp_data_35; ifm_data_44<=temp_data_36;
                                end
                            endcase
                        end
                    end
                    26:begin
                        if(w_cnt ==0)begin
                            ifm_data_15<=1;
                            ifm_data_30<=1;
                            ifm_data_16<=temp_data_0; ifm_data_17<=temp_data_1;  ifm_data_18<=temp_data_2;  ifm_data_19<=temp_data_3;  ifm_data_20<=temp_data_4;  ifm_data_21<=temp_data_5;  ifm_data_22<=temp_data_6;  ifm_data_23<=temp_data_7; ifm_data_24<=temp_data_8; ifm_data_25<=temp_data_9; ifm_data_26<=temp_data_10; ifm_data_27<=temp_data_11; ifm_data_28<=temp_data_12; ifm_data_29<=temp_data_13;
                            ifm_data_31<=temp_data_18; ifm_data_32<=temp_data_19;  ifm_data_33<=temp_data_20;  ifm_data_34<=temp_data_21;  ifm_data_35<=temp_data_22;  ifm_data_36<=temp_data_23;  ifm_data_37<=temp_data_24;  ifm_data_38<=temp_data_25; ifm_data_39<=temp_data_26; ifm_data_40<=temp_data_27; ifm_data_41<=temp_data_28; ifm_data_42<=temp_data_29; ifm_data_43<=temp_data_30; ifm_data_44<=temp_data_31;
                        end else begin
                            ifm_data_29<=1;
                            ifm_data_44<=1;
                            ifm_data_15<=temp_data_0;  ifm_data_16<=temp_data_1; ifm_data_17<=temp_data_2;  ifm_data_18<=temp_data_3;  ifm_data_19<=temp_data_4;  ifm_data_20<=temp_data_5;  ifm_data_21<=temp_data_6;  ifm_data_22<=temp_data_7;  ifm_data_23<=temp_data_8; ifm_data_24<=temp_data_9; ifm_data_25<=temp_data_10; ifm_data_26<=temp_data_11; ifm_data_27<=temp_data_12; ifm_data_28<=temp_data_13;
                            ifm_data_30<=temp_data_18;  ifm_data_31<=temp_data_19; ifm_data_32<=temp_data_20;  ifm_data_33<=temp_data_21;  ifm_data_34<=temp_data_22;  ifm_data_35<=temp_data_23;  ifm_data_36<=temp_data_24;  ifm_data_37<=temp_data_25;  ifm_data_38<=temp_data_26; ifm_data_39<=temp_data_27; ifm_data_40<=temp_data_28; ifm_data_41<=temp_data_29; ifm_data_42<=temp_data_30; ifm_data_43<=temp_data_31;
                        end
                    end
                    13:begin
                        ifm_data_15<=1;
                        ifm_data_30<=1;
                        ifm_data_29<=1;
                        ifm_data_44<=1;
                        case(remain_13)
                            0:begin
                                ifm_data_16<=temp_data_3; ifm_data_17<=temp_data_4;  ifm_data_18<=temp_data_5;  ifm_data_19<=temp_data_6;  ifm_data_20<=temp_data_7;  ifm_data_21<=temp_data_8;  ifm_data_22<=temp_data_9;  ifm_data_23<=temp_data_10; ifm_data_24<=temp_data_11; ifm_data_25<=temp_data_12; ifm_data_26<=temp_data_13; ifm_data_27<=temp_data_14; ifm_data_28<=temp_data_15;
                                ifm_data_31<=temp_data_16; ifm_data_32<=temp_data_17;  ifm_data_33<=temp_data_18;  ifm_data_34<=temp_data_19;  ifm_data_35<=temp_data_20;  ifm_data_36<=temp_data_21;  ifm_data_37<=temp_data_22;  ifm_data_38<=temp_data_23; ifm_data_39<=temp_data_24; ifm_data_40<=temp_data_25; ifm_data_41<=temp_data_26; ifm_data_42<=temp_data_27; ifm_data_43<=temp_data_28;
                            end
                            1:begin
                                ifm_data_16<=temp_data_2; ifm_data_17<=temp_data_3;  ifm_data_18<=temp_data_4;  ifm_data_19<=temp_data_5;  ifm_data_20<=temp_data_6;  ifm_data_21<=temp_data_7;  ifm_data_22<=temp_data_8;  ifm_data_23<=temp_data_9; ifm_data_24<=temp_data_10; ifm_data_25<=temp_data_11; ifm_data_26<=temp_data_12; ifm_data_27<=temp_data_13; ifm_data_28<=temp_data_14;
                                ifm_data_31<=temp_data_19; ifm_data_32<=temp_data_20;  ifm_data_33<=temp_data_21;  ifm_data_34<=temp_data_22;  ifm_data_35<=temp_data_23;  ifm_data_36<=temp_data_24;  ifm_data_37<=temp_data_25;  ifm_data_38<=temp_data_26; ifm_data_39<=temp_data_27; ifm_data_40<=temp_data_28; ifm_data_41<=temp_data_29; ifm_data_42<=temp_data_30; ifm_data_43<=temp_data_31;
                            end
                            2:begin
                                ifm_data_16<=temp_data_1; ifm_data_17<=temp_data_2;  ifm_data_18<=temp_data_3;  ifm_data_19<=temp_data_4;  ifm_data_20<=temp_data_5;  ifm_data_21<=temp_data_6;  ifm_data_22<=temp_data_7;  ifm_data_23<=temp_data_8; ifm_data_24<=temp_data_9; ifm_data_25<=temp_data_10; ifm_data_26<=temp_data_11; ifm_data_27<=temp_data_12; ifm_data_28<=temp_data_13;
                                ifm_data_31<=temp_data_18; ifm_data_32<=temp_data_19;  ifm_data_33<=temp_data_20;  ifm_data_34<=temp_data_21;  ifm_data_35<=temp_data_22;  ifm_data_36<=temp_data_23;  ifm_data_37<=temp_data_24;  ifm_data_38<=temp_data_25; ifm_data_39<=temp_data_26; ifm_data_40<=temp_data_27; ifm_data_41<=temp_data_28; ifm_data_42<=temp_data_29; ifm_data_43<=temp_data_30;
                            end
                            3:begin
                                ifm_data_16<=temp_data_0; ifm_data_17<=temp_data_1;  ifm_data_18<=temp_data_2;  ifm_data_19<=temp_data_3;  ifm_data_20<=temp_data_4;  ifm_data_21<=temp_data_5;  ifm_data_22<=temp_data_6;  ifm_data_23<=temp_data_7; ifm_data_24<=temp_data_8; ifm_data_25<=temp_data_9; ifm_data_26<=temp_data_10; ifm_data_27<=temp_data_11; ifm_data_28<=temp_data_12;
                                ifm_data_31<=temp_data_17; ifm_data_32<=temp_data_18;  ifm_data_33<=temp_data_19;  ifm_data_34<=temp_data_20;  ifm_data_35<=temp_data_21;  ifm_data_36<=temp_data_22;  ifm_data_37<=temp_data_23;  ifm_data_38<=temp_data_24; ifm_data_39<=temp_data_25; ifm_data_40<=temp_data_26; ifm_data_41<=temp_data_27; ifm_data_42<=temp_data_28; ifm_data_43<=temp_data_29;
                            end
                        endcase       
                    end
                endcase
            end else if(buf_conv3_rowlast& bram_hs)begin
                ifm_data_30<=1;  ifm_data_31<=1; ifm_data_32<=1;  ifm_data_33<=1;  ifm_data_34<=1;  ifm_data_35<=1;  ifm_data_36<=1;  ifm_data_37<=1;  ifm_data_38<=1; ifm_data_39<=1; ifm_data_40<=1; ifm_data_41<=1; ifm_data_42<=1; ifm_data_43<=1; ifm_data_44<=1;
                if(read_flag)begin
                    ifm_data_0<=reuse_data_2ifm0[0][15:0]; ifm_data_1<={reuse_data_2ifm0[1][7:0],reuse_data_2ifm0[0][23:16]}; ifm_data_2<=reuse_data_2ifm0[1][23:8];  ifm_data_3<=reuse_data_2ifm0[2][15:0];  ifm_data_4<={reuse_data_2ifm0[3][7:0],reuse_data_2ifm0[2][23:16]};  ifm_data_5<=reuse_data_2ifm0[3][23:8];  ifm_data_6<=reuse_data_2ifm0[4][15:0];  ifm_data_7<={reuse_data_2ifm0[5][7:0],reuse_data_2ifm0[4][23:16]};  ifm_data_8<=reuse_data_2ifm0[5][23:8]; ifm_data_9<=reuse_data_2ifm0[6][15:0]; ifm_data_10<={reuse_data_2ifm0[7][7:0],reuse_data_2ifm0[6][23:16]}; ifm_data_11<=reuse_data_2ifm0[7][23:8]; ifm_data_12<=reuse_data_2ifm0[8][15:0]; ifm_data_13<={reuse_data_2ifm0[9][7:0],reuse_data_2ifm0[8][23:16]}; ifm_data_14<=reuse_data_2ifm0[9][23:8];
                    ifm_data_15<=reuse_data_2ifm0[10][15:0];  ifm_data_16<={reuse_data_2ifm0[11][7:0],reuse_data_2ifm0[10][23:16]}; ifm_data_17<=reuse_data_2ifm0[11][23:8];  ifm_data_18<=reuse_data_2ifm0[12][15:0];  ifm_data_19<={reuse_data_2ifm0[13][7:0],reuse_data_2ifm0[12][23:16]};  ifm_data_20<=reuse_data_2ifm0[13][23:8];  ifm_data_21<=reuse_data_2ifm0[14][15:0];  ifm_data_22<={reuse_data_2ifm0[15][7:0],reuse_data_2ifm0[14][23:16]};  ifm_data_23<=reuse_data_2ifm0[15][23:8]; ifm_data_24<=reuse_data_2ifm0[16][15:0]; ifm_data_25<={reuse_data_2ifm0[17][7:0],reuse_data_2ifm0[16][23:16]}; ifm_data_26<=reuse_data_2ifm0[17][23:8]; ifm_data_27<=reuse_data_2ifm0[18][15:0]; ifm_data_28<={reuse_data_2ifm0[19][7:0],reuse_data_2ifm0[18][23:16]}; ifm_data_29<=reuse_data_2ifm0[19][23:8];
                end else begin
                    ifm_data_0<=reuse_data_2ifm1[0][15:0]; ifm_data_1<={reuse_data_2ifm1[1][7:0],reuse_data_2ifm1[0][23:16]}; ifm_data_2<=reuse_data_2ifm1[1][23:8];  ifm_data_3<=reuse_data_2ifm1[2][15:0];  ifm_data_4<={reuse_data_2ifm1[3][7:0],reuse_data_2ifm1[2][23:16]};  ifm_data_5<=reuse_data_2ifm1[3][23:8];  ifm_data_6<=reuse_data_2ifm1[4][15:0];  ifm_data_7<={reuse_data_2ifm1[5][7:0],reuse_data_2ifm1[4][23:16]};  ifm_data_8<=reuse_data_2ifm1[5][23:8]; ifm_data_9<=reuse_data_2ifm1[6][15:0]; ifm_data_10<={reuse_data_2ifm1[7][7:0],reuse_data_2ifm1[6][23:16]}; ifm_data_11<=reuse_data_2ifm1[7][23:8]; ifm_data_12<=reuse_data_2ifm1[8][15:0]; ifm_data_13<={reuse_data_2ifm1[9][7:0],reuse_data_2ifm1[8][23:16]}; ifm_data_14<=reuse_data_2ifm1[9][23:8];
                    ifm_data_15<=reuse_data_2ifm1[10][15:0];  ifm_data_16<={reuse_data_2ifm1[11][7:0],reuse_data_2ifm1[10][23:16]}; ifm_data_17<=reuse_data_2ifm1[11][23:8];  ifm_data_18<=reuse_data_2ifm1[12][15:0];  ifm_data_19<={reuse_data_2ifm1[13][7:0],reuse_data_2ifm1[12][23:16]};  ifm_data_20<=reuse_data_2ifm1[13][23:8];  ifm_data_21<=reuse_data_2ifm1[14][15:0];  ifm_data_22<={reuse_data_2ifm1[15][7:0],reuse_data_2ifm1[14][23:16]};  ifm_data_23<=reuse_data_2ifm1[15][23:8]; ifm_data_24<=reuse_data_2ifm1[16][15:0]; ifm_data_25<={reuse_data_2ifm1[17][7:0],reuse_data_2ifm1[16][23:16]}; ifm_data_26<=reuse_data_2ifm1[17][23:8]; ifm_data_27<=reuse_data_2ifm1[18][15:0]; ifm_data_28<={reuse_data_2ifm1[19][7:0],reuse_data_2ifm1[18][23:16]}; ifm_data_29<=reuse_data_2ifm1[19][23:8];
                end
            end else if(temp_hs) begin
                if(read_flag)begin
                    ifm_data_0<=reuse_data_2ifm0[0][15:0]; ifm_data_1<={reuse_data_2ifm0[1][7:0],reuse_data_2ifm0[0][23:16]}; ifm_data_2<=reuse_data_2ifm0[1][23:8];  ifm_data_3<=reuse_data_2ifm0[2][15:0];  ifm_data_4<={reuse_data_2ifm0[3][7:0],reuse_data_2ifm0[2][23:16]};  ifm_data_5<=reuse_data_2ifm0[3][23:8];  ifm_data_6<=reuse_data_2ifm0[4][15:0];  ifm_data_7<={reuse_data_2ifm0[5][7:0],reuse_data_2ifm0[4][23:16]};  ifm_data_8<=reuse_data_2ifm0[5][23:8]; ifm_data_9<=reuse_data_2ifm0[6][15:0]; ifm_data_10<={reuse_data_2ifm0[7][7:0],reuse_data_2ifm0[6][23:16]}; ifm_data_11<=reuse_data_2ifm0[7][23:8]; ifm_data_12<=reuse_data_2ifm0[8][15:0]; ifm_data_13<={reuse_data_2ifm0[9][7:0],reuse_data_2ifm0[8][23:16]}; ifm_data_14<=reuse_data_2ifm0[9][23:8];
                    ifm_data_15<=reuse_data_2ifm0[10][15:0];  ifm_data_16<={reuse_data_2ifm0[11][7:0],reuse_data_2ifm0[10][23:16]}; ifm_data_17<=reuse_data_2ifm0[11][23:8];  ifm_data_18<=reuse_data_2ifm0[12][15:0];  ifm_data_19<={reuse_data_2ifm0[13][7:0],reuse_data_2ifm0[12][23:16]};  ifm_data_20<=reuse_data_2ifm0[13][23:8];  ifm_data_21<=reuse_data_2ifm0[14][15:0];  ifm_data_22<={reuse_data_2ifm0[15][7:0],reuse_data_2ifm0[14][23:16]};  ifm_data_23<=reuse_data_2ifm0[15][23:8]; ifm_data_24<=reuse_data_2ifm0[16][15:0]; ifm_data_25<={reuse_data_2ifm0[17][7:0],reuse_data_2ifm0[16][23:16]}; ifm_data_26<=reuse_data_2ifm0[17][23:8]; ifm_data_27<=reuse_data_2ifm0[18][15:0]; ifm_data_28<={reuse_data_2ifm0[19][7:0],reuse_data_2ifm0[18][23:16]}; ifm_data_29<=reuse_data_2ifm0[19][23:8];
                end else begin
                    ifm_data_0<=reuse_data_2ifm1[0][15:0]; ifm_data_1<={reuse_data_2ifm1[1][7:0],reuse_data_2ifm1[0][23:16]}; ifm_data_2<=reuse_data_2ifm1[1][23:8];  ifm_data_3<=reuse_data_2ifm1[2][15:0];  ifm_data_4<={reuse_data_2ifm1[3][7:0],reuse_data_2ifm1[2][23:16]};  ifm_data_5<=reuse_data_2ifm1[3][23:8];  ifm_data_6<=reuse_data_2ifm1[4][15:0];  ifm_data_7<={reuse_data_2ifm1[5][7:0],reuse_data_2ifm1[4][23:16]};  ifm_data_8<=reuse_data_2ifm1[5][23:8]; ifm_data_9<=reuse_data_2ifm1[6][15:0]; ifm_data_10<={reuse_data_2ifm1[7][7:0],reuse_data_2ifm1[6][23:16]}; ifm_data_11<=reuse_data_2ifm1[7][23:8]; ifm_data_12<=reuse_data_2ifm1[8][15:0]; ifm_data_13<={reuse_data_2ifm1[9][7:0],reuse_data_2ifm1[8][23:16]}; ifm_data_14<=reuse_data_2ifm1[9][23:8];
                    ifm_data_15<=reuse_data_2ifm1[10][15:0];  ifm_data_16<={reuse_data_2ifm1[11][7:0],reuse_data_2ifm1[10][23:16]}; ifm_data_17<=reuse_data_2ifm1[11][23:8];  ifm_data_18<=reuse_data_2ifm1[12][15:0];  ifm_data_19<={reuse_data_2ifm1[13][7:0],reuse_data_2ifm1[12][23:16]};  ifm_data_20<=reuse_data_2ifm1[13][23:8];  ifm_data_21<=reuse_data_2ifm1[14][15:0];  ifm_data_22<={reuse_data_2ifm1[15][7:0],reuse_data_2ifm1[14][23:16]};  ifm_data_23<=reuse_data_2ifm1[15][23:8]; ifm_data_24<=reuse_data_2ifm1[16][15:0]; ifm_data_25<={reuse_data_2ifm1[17][7:0],reuse_data_2ifm1[16][23:16]}; ifm_data_26<=reuse_data_2ifm1[17][23:8]; ifm_data_27<=reuse_data_2ifm1[18][15:0]; ifm_data_28<={reuse_data_2ifm1[19][7:0],reuse_data_2ifm1[18][23:16]}; ifm_data_29<=reuse_data_2ifm1[19][23:8];
                end
                case(ifm_width)
                    default:begin
                        if(w_cnt ==0)begin
                            ifm_data_30<=1;
                            case(remain)
                                0:begin ifm_data_31<=temp_data_2; ifm_data_32<=temp_data_3;  ifm_data_33<=temp_data_4;  ifm_data_34<=temp_data_5;  ifm_data_35<=temp_data_6;  ifm_data_36<=temp_data_7;  ifm_data_37<=temp_data_8;  ifm_data_38<=temp_data_9; ifm_data_39<=temp_data_10; ifm_data_40<=temp_data_11; ifm_data_41<=temp_data_12; ifm_data_42<=temp_data_13; ifm_data_43<=temp_data_14; ifm_data_44<=temp_data_15; end
                                2:begin ifm_data_31<=temp_data_0; ifm_data_32<=temp_data_1;  ifm_data_33<=temp_data_2;  ifm_data_34<=temp_data_3;  ifm_data_35<=temp_data_4;  ifm_data_36<=temp_data_5;  ifm_data_37<=temp_data_6;  ifm_data_38<=temp_data_7; ifm_data_39<=temp_data_8; ifm_data_40<=temp_data_9; ifm_data_41<=temp_data_10; ifm_data_42<=temp_data_11; ifm_data_43<=temp_data_12; ifm_data_44<=temp_data_13; end
                            endcase
                        end else if(w_cnt == w_finish_cnt)begin
                            ifm_data_44 <=1;
                            case(remain)
                                0:begin ifm_data_30<=temp_data_2;  ifm_data_31<=temp_data_3; ifm_data_32<=temp_data_4;  ifm_data_33<=temp_data_5;  ifm_data_34<=temp_data_6;  ifm_data_35<=temp_data_7;  ifm_data_36<=temp_data_8;  ifm_data_37<=temp_data_9;  ifm_data_38<=temp_data_10; ifm_data_39<=temp_data_11; ifm_data_40<=temp_data_12; ifm_data_41<=temp_data_13; ifm_data_42<=temp_data_14; ifm_data_43<=temp_data_15; end
                                2:begin ifm_data_30<=temp_data_0;  ifm_data_31<=temp_data_1; ifm_data_32<=temp_data_2;  ifm_data_33<=temp_data_3;  ifm_data_34<=temp_data_4;  ifm_data_35<=temp_data_5;  ifm_data_36<=temp_data_6;  ifm_data_37<=temp_data_7;  ifm_data_38<=temp_data_8; ifm_data_39<=temp_data_9; ifm_data_40<=temp_data_10; ifm_data_41<=temp_data_11; ifm_data_42<=temp_data_12; ifm_data_43<=temp_data_13; end
                            endcase
                        end else begin
                            case(remain)
                                0:begin ifm_data_30<=temp_data_1;  ifm_data_31<=temp_data_2; ifm_data_32<=temp_data_3;  ifm_data_33<=temp_data_4;  ifm_data_34<=temp_data_5;  ifm_data_35<=temp_data_6;  ifm_data_36<=temp_data_7;  ifm_data_37<=temp_data_8;  ifm_data_38<=temp_data_9; ifm_data_39<=temp_data_10; ifm_data_40<=temp_data_11; ifm_data_41<=temp_data_12; ifm_data_42<=temp_data_13; ifm_data_43<=temp_data_14; ifm_data_44<=temp_data_15;end
                                1:begin ifm_data_30<=temp_data_0;  ifm_data_31<=temp_data_1; ifm_data_32<=temp_data_2;  ifm_data_33<=temp_data_3;  ifm_data_34<=temp_data_4;  ifm_data_35<=temp_data_5;  ifm_data_36<=temp_data_6;  ifm_data_37<=temp_data_7;  ifm_data_38<=temp_data_8; ifm_data_39<=temp_data_9; ifm_data_40<=temp_data_10; ifm_data_41<=temp_data_11; ifm_data_42<=temp_data_12; ifm_data_43<=temp_data_13; ifm_data_44<=temp_data_14;end
                                2:begin ifm_data_30<=temp_data_3;  ifm_data_31<=temp_data_4; ifm_data_32<=temp_data_5;  ifm_data_33<=temp_data_6;  ifm_data_34<=temp_data_7;  ifm_data_35<=temp_data_8;  ifm_data_36<=temp_data_9;  ifm_data_37<=temp_data_10;  ifm_data_38<=temp_data_11; ifm_data_39<=temp_data_12; ifm_data_40<=temp_data_13; ifm_data_41<=temp_data_14; ifm_data_42<=temp_data_15; ifm_data_43<=temp_data_16; ifm_data_44<=temp_data_17;end
                                3:begin ifm_data_30<=temp_data_2;  ifm_data_31<=temp_data_3; ifm_data_32<=temp_data_4;  ifm_data_33<=temp_data_5;  ifm_data_34<=temp_data_6;  ifm_data_35<=temp_data_7;  ifm_data_36<=temp_data_8;  ifm_data_37<=temp_data_9;  ifm_data_38<=temp_data_10; ifm_data_39<=temp_data_11; ifm_data_40<=temp_data_12; ifm_data_41<=temp_data_13; ifm_data_42<=temp_data_14; ifm_data_43<=temp_data_15; ifm_data_44<=temp_data_16;end
                            endcase
                        end
                    end
                    13:begin
                        case(remain_13)
                            0: begin ifm_data_30<=1;  ifm_data_31<=temp_data_3; ifm_data_32<=temp_data_4;  ifm_data_33<=temp_data_5;  ifm_data_34<=temp_data_6;  ifm_data_35<=temp_data_7;  ifm_data_36<=temp_data_8;  ifm_data_37<=temp_data_9;  ifm_data_38<=temp_data_10; ifm_data_39<=temp_data_11; ifm_data_40<=temp_data_12; ifm_data_41<=temp_data_13; ifm_data_42<=temp_data_14; ifm_data_43<=temp_data_15; ifm_data_44<=1; end
                            1: begin ifm_data_30<=1;  ifm_data_31<=temp_data_2; ifm_data_32<=temp_data_3;  ifm_data_33<=temp_data_4;  ifm_data_34<=temp_data_5;  ifm_data_35<=temp_data_6;  ifm_data_36<=temp_data_7;  ifm_data_37<=temp_data_8;  ifm_data_38<=temp_data_9; ifm_data_39<=temp_data_10; ifm_data_40<=temp_data_11; ifm_data_41<=temp_data_12; ifm_data_42<=temp_data_13; ifm_data_43<=temp_data_14; ifm_data_44<=1; end
                            2: begin ifm_data_30<=1;  ifm_data_31<=temp_data_1; ifm_data_32<=temp_data_2;  ifm_data_33<=temp_data_3;  ifm_data_34<=temp_data_4;  ifm_data_35<=temp_data_5;  ifm_data_36<=temp_data_6;  ifm_data_37<=temp_data_7;  ifm_data_38<=temp_data_8; ifm_data_39<=temp_data_9; ifm_data_40<=temp_data_10; ifm_data_41<=temp_data_11; ifm_data_42<=temp_data_12; ifm_data_43<=temp_data_13; ifm_data_44<=1; end
                            3: begin ifm_data_30<=1;  ifm_data_31<=temp_data_0; ifm_data_32<=temp_data_1;  ifm_data_33<=temp_data_2;  ifm_data_34<=temp_data_3;  ifm_data_35<=temp_data_4;  ifm_data_36<=temp_data_5;  ifm_data_37<=temp_data_6;  ifm_data_38<=temp_data_7; ifm_data_39<=temp_data_8; ifm_data_40<=temp_data_9; ifm_data_41<=temp_data_10; ifm_data_42<=temp_data_11; ifm_data_43<=temp_data_12; ifm_data_44<=1; end
                        endcase
                    end
                endcase
            end
        end
    end
    
endmodule



/*
            ifm_data_0<=temp_data_ ; ifm_data_1<=temp_data_; ifm_data_2<=temp_data_;  ifm_data_3<=temp_data_;  ifm_data_4<=temp_data_;  ifm_data_5<=temp_data_;  ifm_data_6<=temp_data_;  ifm_data_7<=temp_data_;  ifm_data_8<=temp_data_; ifm_data_9<=temp_data_; ,ifm_data_10<=temp_data_; ifm_data_11<=temp_data_; ifm_data_12<=temp_data_; ifm_data_13<=temp_data_; ifm_data_14<=temp_data_;
            ifm_data_15<=temp_data_;  ifm_data_16<=temp_data_; ifm_data_17<=temp_data_;  ifm_data_18<=temp_data_;  ifm_data_19<=temp_data_;  ifm_data_20<=temp_data_;  ifm_data_21<=temp_data_;  ifm_data_22<=temp_data_;  ifm_data_23<=temp_data_; ifm_data_24<=temp_data_; ifm_data_25<=temp_data_; ifm_data_26<=temp_data_; ifm_data_27<=temp_data_; ifm_data_28<=temp_data_; ifm_data_29<=temp_data_;
            ifm_data_30<=temp_data_;  ifm_data_31<=temp_data_; ifm_data_32<=temp_data_;  ifm_data_33<=temp_data_;  ifm_data_34<=temp_data_;  ifm_data_35<=temp_data_;  ifm_data_36<=temp_data_;  ifm_data_37<=temp_data_;  ifm_data_38<=temp_data_; ifm_data_39<=temp_data_; ifm_data_40<=temp_data_; ifm_data_41<=temp_data_; ifm_data_42<=temp_data_; ifm_data_43<=temp_data_; ifm_data_44<=temp_data_;
*/
